`ifndef VERIF_COMPONENTS_SVH
`define VERIF_COMPONENTS_SVH

    `include "components/transaction_base.svh"
    `include "components/sequence_base.svh"
    `include "components/host_guest_channel.svh"
    `include "components/driver_base.svh"
    `include "components/scoreboard_base.svh"
    `include "components/monitor_base.svh"
    `include "components/env_base.svh"
    `include "components/test_config_base.svh"

`endif  // VERIF_COMPONENTS_SVH

