package uart_tests_pkg;

    import uart_tb_pkg::*;
    import axi4l_pkg::*;

`include "uart_test_base.sv"
`include "uart_test_scratch.sv"

endpackage: uart_tests_pkg
