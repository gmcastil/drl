virtual class test_base extends component_base;

    function new(string name = "test_base", component_base parent = null);
        super.new(name, parent);
    endfunction: new

endclass: test_base

