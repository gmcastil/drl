package common_pkg;

`include "data_types.sv"

    // Global default log level (can be overridden)
    localparam  log_level_t     DEFAULT_LOG_LEVEL = LOG_INFO;

endpackage: common_pkg
