package base_pkg;

    import common_pkg::*;

`include "logger.sv"
`include "object_base.sv"

`include "component_base.sv"
`include "config_db.sv"
`include "transaction_base.sv"
`include "sequence_base.sv"
`include "sequencer_base.sv"
`include "driver_base.sv"
`include "env_base.sv"
`include "monitor_base.sv"
`include "scoreboard_base.sv"
`include "test_base.sv"

endpackage: base_pkg

