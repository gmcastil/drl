virtual class monitor_base extends component_base;

    function new(string name, component_base parent);
        super.new(name, parent);
    endfunction: new

endclass: monitor_base
