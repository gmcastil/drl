class test_config_base extends object_base;

    function new(string name);
        super.new(name);
    endfunction: new

endclass: test_config_base

