`ifndef VERIF_PKG_SVH
`define VERIF_PKG_SVH

`include "verif_macros.svh"

package verif_pkg;

    `include "types/verif_types.svh"
    `include "base/verif_base.svh"
    `include "components/verif_components.svh"

endpackage: verif_pkg

`endif  // VERIF_PKG_SVH

