`ifndef VERIF_MACROS_SVH
`define VERIF_MACROS_SVH

`include "macros/verif_logging.svh"

`endif  // VERIF_MACROS_SVH

