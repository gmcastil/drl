virtual class sequence_base extends object_base;

    function new(string name);
        super.new(name);
    endfunction;

endclass: sequence_base
