package uart_tests_pkg;

    import uart_tb_pkg::*;

`include "uart_test_base.sv"

endpackage: uart_tests_pkg
