virtual class env_base extends component_base;

    function new(string name = "env_base", component_base parent = null);
        super.new(name, parent);
    endfunction: new

endclass: env_base

