`ifndef VERIF_TYPES_SVH
`define VERIF_TYPES_SVH

    `include "types/logging_types.svh"

`endif  // VERIF_TYPES_SVH

