package common_pkg;

`include "data_types.sv"
`include "macros.svh"

endpackage: common_pkg
