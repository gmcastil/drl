package uart_tb_pkg;

    import axi4l_pkg::*;

`include "uart_config.sv"
`include "uart_sequencer.sv"
`include "uart_env.sv"

endpackage: uart_tb_pkg

