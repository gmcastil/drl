package tests_pkg;

    import common_pkg::*;
    import base_pkg::*;

`include "base_test.sv"
`include "env_test.sv"

endpackage: tests_pkg

