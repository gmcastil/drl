`ifndef VERIF_BASE_SVH
`define VERIF_BASE_SVH

    typedef class logger;

    `include "base/object_base.svh"
    `include "base/component_base.svh"
    `include "base/config_db.svh"
    `include "base/logger.svh"
    `include "base/objection_mgr.svh"
    `include "base/test_case_base.svh"
    `include "base/test_factory.svh"
    `include "base/test_root.svh"

`endif  // VERIF_BASE_SVH

